use std.textio.all;entity a is end;architecture b of a is
begin write(output,"10\n11\n12\n13\n14\n15\n16\n17\n20\n22\n24\n31\n100\n121\n10000");end;