use std.textio.all;entity a is end;architecture b of a is
begin write(output,"v");end;