entity e is end;architecture a of e is
begin
process
begin
while 1>0 loop end loop;end process;end;